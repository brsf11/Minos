`timescale 1ns/1ps
module testbench();

    reg CLK,rst_n;
    reg[31:0] ROMData,RAMData;
    wire[31:0] IFPC,RADDR,WADDR,WData;
    wire[1:0] RWHBS,WWHBS;
    wire WE;

    RISCVCore riscvcore(
        .CLK(CLK),
        .rst_n(rst_n),
        .ROMData(ROMData),
        .RAMData(RAMData),
        .IFPC(IFPC),
        .RADDR(RADDR),
        .WADDR(WADDR),
        .WData(WData),
        .RWHBS(RWHBS),
        .WWHBS(WWHBS),
        .WE(WE)
    );


    initial begin
        rst_n=0;
        #10;
        rst_n=1;
        ROMData=32'h0c848493;
        #10;
        ROMData=32'h0c848493;
        #10;
        ROMData=32'h0c848493;
        #10;
        ROMData=32'h0c848493;
        #10;
        ROMData=32'h0c848493;
        #10;
        ROMData=32'h0c848493;
        #10;
        ROMData=32'h0c848493;
        #10;
        ROMData=32'h0c848493;
        #10;
        ROMData=32'h0c848493;
        #10;
        ROMData=32'h0c848493;
        #10;
        ROMData=32'h0c848493;
        #10;
        ROMData=32'h0c848493;
        #10;
        
        
    end

    initial begin
        $dumpfile("wave.vcd");
        $dumpvars(0,testbench);
    end

    initial begin
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
    end

endmodule