`timescale 1ns/1ps
module testbench();

    reg CLK,rst_n;

    top top(
        .CLK(CLK),
        .rst_n(rst_n)
    );

    initial begin
        rst_n=0;
        #10;
        rst_n=1;
    end

    initial begin
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
        CLK=0;
        #5;
        CLK=1;
        #5;
    end

    initial begin
        $dumpfile("wave.vcd");
        $dumpvars(0,testbench);
    end 

endmodule